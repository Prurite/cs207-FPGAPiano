`define nNU  9'b00_0000000

`define nC3  9'b10_0000001
`define nD3  9'b10_0000010
`define nE3  9'b10_0000100
`define nF3  9'b10_0001000
`define nG3  9'b10_0010000
`define nA3  9'b10_0100000
`define nB3  9'b10_1000000

`define nC4  9'b00_0000001
`define nD4  9'b00_0000010
`define nE4  9'b00_0000100
`define nF4  9'b00_0001000
`define nG4  9'b00_0010000
`define nA4  9'b00_0100000
`define nB4  9'b00_1000000

`define nC5  9'b01_0000001
`define nD5  9'b01_0000010
`define nE5  9'b01_0000100
`define nF5  9'b01_0001000
`define nG5  9'b01_0010000
`define nA5  9'b01_0100000
`define nB5  9'b01_1000000