module pageMainMenu(
    input clk,
    input rst,
	input UserInput user_in,
    output ProgramOutput prog_out
);
endmodule
