/* Original file
 * https://github.com/Derek-X-Wang/VGA-Text-Generator/blob/master/VGA-Text-Generator.srcs/sources_1/new/Font_Rom.vhd
 * Rewritten in SystemVerilog
 */

module Font_Rom (
    input logic clk,
    input integer addr,
    output logic [7:0] fontRow
);

    // Parameters for font dimensions
    parameter integer FONT_WIDTH = 8;
    parameter integer CHARACTERS = 128;
    parameter integer ROWS_PER_CHAR = 16;
    parameter integer ROM_SIZE = 2048; // 2^11

    // Define ROM type
    typedef logic [FONT_WIDTH-1:0] rom_row_t;
    typedef rom_row_t rom_t [ROM_SIZE];

    // ROM initialization with font data
    rom_t ROM = {
        // NUL: code x00
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // SOH: code x01
        8'b00000000,
        8'b00000000,
        8'b01111110,
        8'b10000001,
        8'b10100101,
        8'b10000001,
        8'b10000001,
        8'b10111101,
        8'b10011001,
        8'b10000001,
        8'b10000001,
        8'b01111110,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // STX: code x02
        8'b00000000,
        8'b00000000,
        8'b01111110,
        8'b11111111,
        8'b11011011,
        8'b11111111,
        8'b11111111,
        8'b11000011,
        8'b11100111,
        8'b11111111,
        8'b11111111,
        8'b01111110,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // ETX: code x03
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b01101100,
        8'b11111110,
        8'b11111110,
        8'b11111110,
        8'b11111110,
        8'b01111100,
        8'b00111000,
        8'b00010000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // EOT: code x04
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00010000,
        8'b00111000,
        8'b01111100,
        8'b11111110,
        8'b01111100,
        8'b00111000,
        8'b00010000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // ENQ: code x05
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00011000,
        8'b00111100,
        8'b00111100,
        8'b11100111,
        8'b11100111,
        8'b11100111,
        8'b00011000,
        8'b00011000,
        8'b00111100,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // ACK: code x06
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00011000,
        8'b00111100,
        8'b01111110,
        8'b11111111,
        8'b11111111,
        8'b01111110,
        8'b00011000,
        8'b00011000,
        8'b00111100,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // BEL: code x07
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00011000,
        8'b00111100,
        8'b00111100,
        8'b00011000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // BS: code x08
        8'b11111111,
        8'b11111111,
        8'b11111111,
        8'b11111111,
        8'b11111111,
        8'b11111111,
        8'b11100111,
        8'b11000011,
        8'b11000011,
        8'b11100111,
        8'b11111111,
        8'b11111111,
        8'b11111111,
        8'b11111111,
        8'b11111111,
        8'b11111111,
        // HT: code x09
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00111100,
        8'b01100110,
        8'b01000010,
        8'b01000010,
        8'b01100110,
        8'b00111100,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // LF: code x0a
        8'b11111111,
        8'b11111111,
        8'b11111111,
        8'b11111111,
        8'b11111111,
        8'b11000011,
        8'b10011001,
        8'b10111101,
        8'b10111101,
        8'b10011001,
        8'b11000011,
        8'b11111111,
        8'b11111111,
        8'b11111111,
        8'b11111111,
        8'b11111111,
        // code x0b
        8'b00000000,
        8'b00000000,
        8'b00011110,
        8'b00001110,
        8'b00011010,
        8'b00110010,
        8'b01111000,
        8'b11001100,
        8'b11001100,
        8'b11001100,
        8'b11001100,
        8'b01111000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x0c
        8'b00000000,
        8'b00000000,
        8'b00111100,
        8'b01100110,
        8'b01100110,
        8'b01100110,
        8'b01100110,
        8'b00111100,
        8'b00011000,
        8'b01111110,
        8'b00011000,
        8'b00011000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x0d
        8'b00000000,
        8'b00000000,
        8'b00111111,
        8'b00110011,
        8'b00111111,
        8'b00110000,
        8'b00110000,
        8'b00110000,
        8'b00110000,
        8'b01110000,
        8'b11110000,
        8'b11100000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x0e
        8'b00000000,
        8'b00000000,
        8'b01111111,
        8'b01100011,
        8'b01111111,
        8'b01100011,
        8'b01100011,
        8'b01100011,
        8'b01100011,
        8'b01100111,
        8'b11100111,
        8'b11100110,
        8'b11000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x0f
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00011000,
        8'b00011000,
        8'b11011011,
        8'b00111100,
        8'b11100111,
        8'b00111100,
        8'b11011011,
        8'b00011000,
        8'b00011000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x10
        8'b00000000,
        8'b10000000,
        8'b11000000,
        8'b11100000,
        8'b11110000,
        8'b11111000,
        8'b11111110,
        8'b11111000,
        8'b11110000,
        8'b11100000,
        8'b11000000,
        8'b10000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x11
        8'b00000000,
        8'b00000010,
        8'b00000110,
        8'b00001110,
        8'b00011110,
        8'b00111110,
        8'b11111110,
        8'b00111110,
        8'b00011110,
        8'b00001110,
        8'b00000110,
        8'b00000010,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x12
        8'b00000000,
        8'b00000000,
        8'b00011000,
        8'b00111100,
        8'b01111110,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b01111110,
        8'b00111100,
        8'b00011000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x13
        8'b00000000,
        8'b00000000,
        8'b01100110,
        8'b01100110,
        8'b01100110,
        8'b01100110,
        8'b01100110,
        8'b01100110,
        8'b01100110,
        8'b00000000,
        8'b01100110,
        8'b01100110,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x14
        8'b00000000,
        8'b00000000,
        8'b01111111,
        8'b11011011,
        8'b11011011,
        8'b11011011,
        8'b01111011,
        8'b00011011,
        8'b00011011,
        8'b00011011,
        8'b00011011,
        8'b00011011,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x15
        8'b00000000,
        8'b01111100,
        8'b11000110,
        8'b01100000,
        8'b00111000,
        8'b01101100,
        8'b11000110,
        8'b11000110,
        8'b01101100,
        8'b00111000,
        8'b00001100,
        8'b11000110,
        8'b01111100,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x16
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b11111110,
        8'b11111110,
        8'b11111110,
        8'b11111110,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x17
        8'b00000000,
        8'b00000000,
        8'b00011000,
        8'b00111100,
        8'b01111110,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b01111110,
        8'b00111100,
        8'b00011000,
        8'b01111110,
        8'b00110000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x18
        8'b00000000,
        8'b00000000,
        8'b00011000,
        8'b00111100,
        8'b01111110,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x19
        8'b00000000,
        8'b00000000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b01111110,
        8'b00111100,
        8'b00011000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x1a
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00011000,
        8'b00001100,
        8'b11111110,
        8'b00001100,
        8'b00011000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x1b
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00110000,
        8'b01100000,
        8'b11111110,
        8'b01100000,
        8'b00110000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x1c
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b11000000,
        8'b11000000,
        8'b11000000,
        8'b11111110,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x1d
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00100100,
        8'b01100110,
        8'b11111111,
        8'b01100110,
        8'b00100100,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x1e
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00010000,
        8'b00111000,
        8'b00111000,
        8'b01111100,
        8'b01111100,
        8'b11111110,
        8'b11111110,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x1f
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b11111110,
        8'b11111110,
        8'b01111100,
        8'b01111100,
        8'b00111000,
        8'b00111000,
        8'b00010000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x20
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x21
        8'b00000000,
        8'b00000000,
        8'b00011000,
        8'b00111100,
        8'b00111100,
        8'b00111100,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00000000,
        8'b00011000,
        8'b00011000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x22
        8'b00000000,
        8'b01100110,
        8'b01100110,
        8'b01100110,
        8'b00100100,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x23
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b01101100,
        8'b01101100,
        8'b11111110,
        8'b01101100,
        8'b01101100,
        8'b01101100,
        8'b11111110,
        8'b01101100,
        8'b01101100,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x24
        8'b00011000,
        8'b00011000,
        8'b01111100,
        8'b11000110,
        8'b11000010,
        8'b11000000,
        8'b01111100,
        8'b00000110,
        8'b00000110,
        8'b10000110,
        8'b11000110,
        8'b01111100,
        8'b00011000,
        8'b00011000,
        8'b00000000,
        8'b00000000,
        // code x25
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b11000010,
        8'b11000110,
        8'b00001100,
        8'b00011000,
        8'b00110000,
        8'b01100000,
        8'b11000110,
        8'b10000110,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x26
        8'b00000000,
        8'b00000000,
        8'b00111000,
        8'b01101100,
        8'b01101100,
        8'b00111000,
        8'b01110110,
        8'b11011100,
        8'b11001100,
        8'b11001100,
        8'b11001100,
        8'b01110110,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x27
        8'b00000000,
        8'b00110000,
        8'b00110000,
        8'b00110000,
        8'b01100000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x28
        8'b00000000,
        8'b00000000,
        8'b00001100,
        8'b00011000,
        8'b00110000,
        8'b00110000,
        8'b00110000,
        8'b00110000,
        8'b00110000,
        8'b00110000,
        8'b00011000,
        8'b00001100,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x29
        8'b00000000,
        8'b00000000,
        8'b00110000,
        8'b00011000,
        8'b00001100,
        8'b00001100,
        8'b00001100,
        8'b00001100,
        8'b00001100,
        8'b00001100,
        8'b00011000,
        8'b00110000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x2a
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b01100110,
        8'b00111100,
        8'b11111111,
        8'b00111100,
        8'b01100110,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x2b
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00011000,
        8'b00011000,
        8'b01111110,
        8'b00011000,
        8'b00011000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x2c
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00110000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x2d
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b01111110,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x2e
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00011000,
        8'b00011000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x2f
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000010,
        8'b00000110,
        8'b00001100,
        8'b00011000,
        8'b00110000,
        8'b01100000,
        8'b11000000,
        8'b10000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // 0: code x30
        8'b00000000,
        8'b00000000,
        8'b01111100,
        8'b11000110,
        8'b11000110,
        8'b11001110,
        8'b11011110,
        8'b11110110,
        8'b11100110,
        8'b11000110,
        8'b11000110,
        8'b01111100,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // 1: code x31
        8'b00000000,
        8'b00000000,
        8'b00011000,
        8'b00111000,
        8'b01111000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b01111110,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // 2: code x32
        8'b00000000,
        8'b00000000,
        8'b01111100,
        8'b11000110,
        8'b00000110,
        8'b00001100,
        8'b00011000,
        8'b00110000,
        8'b01100000,
        8'b11000000,
        8'b11000110,
        8'b11111110,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // 3: code x33
        8'b00000000,
        8'b00000000,
        8'b01111100,
        8'b11000110,
        8'b00000110,
        8'b00000110,
        8'b00111100,
        8'b00000110,
        8'b00000110,
        8'b00000110,
        8'b11000110,
        8'b01111100,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // 4: code x34
        8'b00000000,
        8'b00000000,
        8'b00001100,
        8'b00011100,
        8'b00111100,
        8'b01101100,
        8'b11001100,
        8'b11111110,
        8'b00001100,
        8'b00001100,
        8'b00001100,
        8'b00011110,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x35
        8'b00000000,
        8'b00000000,
        8'b11111110,
        8'b11000000,
        8'b11000000,
        8'b11000000,
        8'b11111100,
        8'b00000110,
        8'b00000110,
        8'b00000110,
        8'b11000110,
        8'b01111100,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x36
        8'b00000000,
        8'b00000000,
        8'b00111000,
        8'b01100000,
        8'b11000000,
        8'b11000000,
        8'b11111100,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b01111100,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x37
        8'b00000000,
        8'b00000000,
        8'b11111110,
        8'b11000110,
        8'b00000110,
        8'b00000110,
        8'b00001100,
        8'b00011000,
        8'b00110000,
        8'b00110000,
        8'b00110000,
        8'b00110000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x38
        8'b00000000,
        8'b00000000,
        8'b01111100,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b01111100,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b01111100,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x39
        8'b00000000,
        8'b00000000,
        8'b01111100,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b01111110,
        8'b00000110,
        8'b00000110,
        8'b00000110,
        8'b00001100,
        8'b01111000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x3a
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00011000,
        8'b00011000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00011000,
        8'b00011000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x3b
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00011000,
        8'b00011000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00011000,
        8'b00011000,
        8'b00110000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x3c
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000110,
        8'b00001100,
        8'b00011000,
        8'b00110000,
        8'b01100000,
        8'b00110000,
        8'b00011000,
        8'b00001100,
        8'b00000110,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x3d
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b01111110,
        8'b00000000,
        8'b00000000,
        8'b01111110,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x3e
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b01100000,
        8'b00110000,
        8'b00011000,
        8'b00001100,
        8'b00000110,
        8'b00001100,
        8'b00011000,
        8'b00110000,
        8'b01100000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x3f
        8'b00000000,
        8'b00000000,
        8'b01111100,
        8'b11000110,
        8'b11000110,
        8'b00001100,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00000000,
        8'b00011000,
        8'b00011000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x40
        8'b00000000,
        8'b00000000,
        8'b01111100,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b11011110,
        8'b11011110,
        8'b11011110,
        8'b11011100,
        8'b11000000,
        8'b01111100,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // A: code x41
        8'b00000000,
        8'b00000000,
        8'b00010000,
        8'b00111000,
        8'b01101100,
        8'b11000110,
        8'b11000110,
        8'b11111110,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // B: code x42
        8'b00000000,
        8'b00000000,
        8'b11111100,
        8'b01100110,
        8'b01100110,
        8'b01100110,
        8'b01111100,
        8'b01100110,
        8'b01100110,
        8'b01100110,
        8'b01100110,
        8'b11111100,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // C: code x43
        8'b00000000,
        8'b00000000,
        8'b00111100,
        8'b01100110,
        8'b11000010,
        8'b11000000,
        8'b11000000,
        8'b11000000,
        8'b11000000,
        8'b11000010,
        8'b01100110,
        8'b00111100,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // D: code x44
        8'b00000000,
        8'b00000000,
        8'b11111000,
        8'b01101100,
        8'b01100110,
        8'b01100110,
        8'b01100110,
        8'b01100110,
        8'b01100110,
        8'b01100110,
        8'b01101100,
        8'b11111000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x45
        8'b00000000,
        8'b00000000,
        8'b11111110,
        8'b01100110,
        8'b01100010,
        8'b01101000,
        8'b01111000,
        8'b01101000,
        8'b01100000,
        8'b01100010,
        8'b01100110,
        8'b11111110,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x46
        8'b00000000,
        8'b00000000,
        8'b11111110,
        8'b01100110,
        8'b01100010,
        8'b01101000,
        8'b01111000,
        8'b01101000,
        8'b01100000,
        8'b01100000,
        8'b01100000,
        8'b11110000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x47
        8'b00000000,
        8'b00000000,
        8'b00111100,
        8'b01100110,
        8'b11000010,
        8'b11000000,
        8'b11000000,
        8'b11011110,
        8'b11000110,
        8'b11000110,
        8'b01100110,
        8'b00111010,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // H: code x48
        8'b00000000,
        8'b00000000,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b11111110,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // I: code x49
        8'b00000000,
        8'b00000000,
        8'b00111100,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00111100,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // J: code x4a
        8'b00000000,
        8'b00000000,
        8'b00011110,
        8'b00001100,
        8'b00001100,
        8'b00001100,
        8'b00001100,
        8'b00001100,
        8'b11001100,
        8'b11001100,
        8'b11001100,
        8'b01111000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // K: code x4b
        8'b00000000,
        8'b00000000,
        8'b11100110,
        8'b01100110,
        8'b01100110,
        8'b01101100,
        8'b01111000,
        8'b01111000,
        8'b01101100,
        8'b01100110,
        8'b01100110,
        8'b11100110,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // L: code x4c
        8'b00000000,
        8'b00000000,
        8'b11110000,
        8'b01100000,
        8'b01100000,
        8'b01100000,
        8'b01100000,
        8'b01100000,
        8'b01100000,
        8'b01100010,
        8'b01100110,
        8'b11111110,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // M: code x4d
        8'b00000000,
        8'b00000000,
        8'b11000011,
        8'b11100111,
        8'b11111111,
        8'b11111111,
        8'b11011011,
        8'b11000011,
        8'b11000011,
        8'b11000011,
        8'b11000011,
        8'b11000011,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // N: code x4e
        8'b00000000,
        8'b00000000,
        8'b11000110,
        8'b11100110,
        8'b11110110,
        8'b11111110,
        8'b11011110,
        8'b11001110,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // O: code x4f
        8'b00000000,
        8'b00000000,
        8'b01111100,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b01111100,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // P: code x50
        8'b00000000,
        8'b00000000,
        8'b11111100,
        8'b01100110,
        8'b01100110,
        8'b01100110,
        8'b01111100,
        8'b01100000,
        8'b01100000,
        8'b01100000,
        8'b01100000,
        8'b11110000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // Q: code x510
        8'b00000000,
        8'b00000000,
        8'b01111100,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b11010110,
        8'b11011110,
        8'b01111100,
        8'b00001100,
        8'b00001110,
        8'b00000000,
        8'b00000000,
        // code x52
        8'b00000000,
        8'b00000000,
        8'b11111100,
        8'b01100110,
        8'b01100110,
        8'b01100110,
        8'b01111100,
        8'b01101100,
        8'b01100110,
        8'b01100110,
        8'b01100110,
        8'b11100110,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x53
        8'b00000000,
        8'b00000000,
        8'b01111100,
        8'b11000110,
        8'b11000110,
        8'b01100000,
        8'b00111000,
        8'b00001100,
        8'b00000110,
        8'b11000110,
        8'b11000110,
        8'b01111100,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x54
        8'b00000000,
        8'b00000000,
        8'b11111111,
        8'b11011011,
        8'b10011001,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00111100,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x55
        8'b00000000,
        8'b00000000,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b01111100,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x56
        8'b00000000,
        8'b00000000,
        8'b11000011,
        8'b11000011,
        8'b11000011,
        8'b11000011,
        8'b11000011,
        8'b11000011,
        8'b11000011,
        8'b01100110,
        8'b00111100,
        8'b00011000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x57
        8'b00000000,
        8'b00000000,
        8'b11000011,
        8'b11000011,
        8'b11000011,
        8'b11000011,
        8'b11000011,
        8'b11011011,
        8'b11011011,
        8'b11111111,
        8'b01100110,
        8'b01100110,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x58
        8'b00000000,
        8'b00000000,
        8'b11000011,
        8'b11000011,
        8'b01100110,
        8'b00111100,
        8'b00011000,
        8'b00011000,
        8'b00111100,
        8'b01100110,
        8'b11000011,
        8'b11000011,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x59
        8'b00000000,
        8'b00000000,
        8'b11000011,
        8'b11000011,
        8'b11000011,
        8'b01100110,
        8'b00111100,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00111100,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x5a
        8'b00000000,
        8'b00000000,
        8'b11111111,
        8'b11000011,
        8'b10000110,
        8'b00001100,
        8'b00011000,
        8'b00110000,
        8'b01100000,
        8'b11000001,
        8'b11000011,
        8'b11111111,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x5b
        8'b00000000,
        8'b00000000,
        8'b00111100,
        8'b00110000,
        8'b00110000,
        8'b00110000,
        8'b00110000,
        8'b00110000,
        8'b00110000,
        8'b00110000,
        8'b00110000,
        8'b00111100,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x5c
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b10000000,
        8'b11000000,
        8'b11100000,
        8'b01110000,
        8'b00111000,
        8'b00011100,
        8'b00001110,
        8'b00000110,
        8'b00000010,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x5d
        8'b00000000,
        8'b00000000,
        8'b00111100,
        8'b00001100,
        8'b00001100,
        8'b00001100,
        8'b00001100,
        8'b00001100,
        8'b00001100,
        8'b00001100,
        8'b00001100,
        8'b00111100,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x5e
        8'b00010000,
        8'b00111000,
        8'b01101100,
        8'b11000110,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x5f
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b11111111,
        8'b00000000,
        8'b00000000,
        // code x60
        8'b00110000,
        8'b00110000,
        8'b00011000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // a: code x61
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b01111000,
        8'b00001100,
        8'b01111100,
        8'b11001100,
        8'b11001100,
        8'b11001100,
        8'b01110110,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // b: code x62
        8'b00000000,
        8'b00000000,
        8'b11100000,
        8'b01100000,
        8'b01100000,
        8'b01111000,
        8'b01101100,
        8'b01100110,
        8'b01100110,
        8'b01100110,
        8'b01100110,
        8'b01111100,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // c: code x63
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b01111100,
        8'b11000110,
        8'b11000000,
        8'b11000000,
        8'b11000000,
        8'b11000110,
        8'b01111100,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // d: code x64
        8'b00000000,
        8'b00000000,
        8'b00011100,
        8'b00001100,
        8'b00001100,
        8'b00111100,
        8'b01101100,
        8'b11001100,
        8'b11001100,
        8'b11001100,
        8'b11001100,
        8'b01110110,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // e: code x65
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b01111100,
        8'b11000110,
        8'b11111110,
        8'b11000000,
        8'b11000000,
        8'b11000110,
        8'b01111100,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // f: code x66
        8'b00000000,
        8'b00000000,
        8'b00111000,
        8'b01101100,
        8'b01100100,
        8'b01100000,
        8'b11110000,
        8'b01100000,
        8'b01100000,
        8'b01100000,
        8'b01100000,
        8'b11110000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // g: code x67
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b01110110,
        8'b11001100,
        8'b11001100,
        8'b11001100,
        8'b11001100,
        8'b11001100,
        8'b01111100,
        8'b00001100,
        8'b11001100,
        8'b01111000,
        8'b00000000,
        // h: code x68
        8'b00000000,
        8'b00000000,
        8'b11100000,
        8'b01100000,
        8'b01100000,
        8'b01101100,
        8'b01110110,
        8'b01100110,
        8'b01100110,
        8'b01100110,
        8'b01100110,
        8'b11100110,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // i: code x69
        8'b00000000,
        8'b00000000,
        8'b00011000,
        8'b00011000,
        8'b00000000,
        8'b00111000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00111100,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // j: code x6a
        8'b00000000,
        8'b00000000,
        8'b00000110,
        8'b00000110,
        8'b00000000,
        8'b00001110,
        8'b00000110,
        8'b00000110,
        8'b00000110,
        8'b00000110,
        8'b00000110,
        8'b00000110,
        8'b01100110,
        8'b01100110,
        8'b00111100,
        8'b00000000,
        // k: code x6b
        8'b00000000,
        8'b00000000,
        8'b11100000,
        8'b01100000,
        8'b01100000,
        8'b01100110,
        8'b01101100,
        8'b01111000,
        8'b01111000,
        8'b01101100,
        8'b01100110,
        8'b11100110,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // l: code x6c
        8'b00000000,
        8'b00000000,
        8'b00111000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00111100,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // m: code x6d
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b11100110,
        8'b11111111,
        8'b11011011,
        8'b11011011,
        8'b11011011,
        8'b11011011,
        8'b11011011,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // n: code x6e
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b11011100,
        8'b01100110,
        8'b01100110,
        8'b01100110,
        8'b01100110,
        8'b01100110,
        8'b01100110,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // o: code x6f
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b01111100,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b01111100,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x70
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b11011100,
        8'b01100110,
        8'b01100110,
        8'b01100110,
        8'b01100110,
        8'b01100110,
        8'b01111100,
        8'b01100000,
        8'b01100000,
        8'b11110000,
        8'b00000000,
        // code x71
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b01110110,
        8'b11001100,
        8'b11001100,
        8'b11001100,
        8'b11001100,
        8'b11001100,
        8'b01111100,
        8'b00001100,
        8'b00001100,
        8'b00011110,
        8'b00000000,
        // code x72
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b11011100,
        8'b01110110,
        8'b01100110,
        8'b01100000,
        8'b01100000,
        8'b01100000,
        8'b11110000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x73
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b01111100,
        8'b11000110,
        8'b01100000,
        8'b00111000,
        8'b00001100,
        8'b11000110,
        8'b01111100,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x74
        8'b00000000,
        8'b00000000,
        8'b00010000,
        8'b00110000,
        8'b00110000,
        8'b11111100,
        8'b00110000,
        8'b00110000,
        8'b00110000,
        8'b00110000,
        8'b00110110,
        8'b00011100,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x75
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b11001100,
        8'b11001100,
        8'b11001100,
        8'b11001100,
        8'b11001100,
        8'b11001100,
        8'b01110110,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x76
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b11000011,
        8'b11000011,
        8'b11000011,
        8'b11000011,
        8'b01100110,
        8'b00111100,
        8'b00011000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x77
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b11000011,
        8'b11000011,
        8'b11000011,
        8'b11011011,
        8'b11011011,
        8'b11111111,
        8'b01100110,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x78
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b11000011,
        8'b01100110,
        8'b00111100,
        8'b00011000,
        8'b00111100,
        8'b01100110,
        8'b11000011,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x79
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b01111110,
        8'b00000110,
        8'b00001100,
        8'b11111000,
        8'b00000000,
        // code x7a
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b11111110,
        8'b11001100,
        8'b00011000,
        8'b00110000,
        8'b01100000,
        8'b11000110,
        8'b11111110,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x7b
        8'b00000000,
        8'b00000000,
        8'b00001110,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b01110000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00001110,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x7c
        8'b00000000,
        8'b00000000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00000000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x7d
        8'b00000000,
        8'b00000000,
        8'b01110000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00001110,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b00011000,
        8'b01110000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x7e
        8'b00000000,
        8'b00000000,
        8'b01110110,
        8'b11011100,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        // code x7f
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00010000,
        8'b00111000,
        8'b01101100,
        8'b11000110,
        8'b11000110,
        8'b11000110,
        8'b11111110,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000,
        8'b00000000
    };

    // Sequential logic to read from ROM
    always_ff @(posedge clk) begin
        fontRow <= ROM[addr];
    end

endmodule
