`include "header.svh"

module pageMenu(
    input logic clk, prog_clk, rst,
    input UserInput user_in,
    output ProgramOutput menu_out,
    output byte read_chart_id,
    input Chart chart_data,
    output logic auto_play
);
    localparam UP = 4'b1000;
    localparam DOWN = 4'b0100;
    localparam LEFT = 4'b0010;
    localparam RIGHT = 4'b0001;
    byte cur_pos;
    byte chart_id;
    ScreenText text;
    SegDisplayText seg;
    TopState state;

    assign menu_out.text = text;
    assign menu_out.seg = seg;
    assign menu_out.state = state;
    
    always @(posedge prog_clk) begin
        if (rst) begin
            auto_play <= 0;
            cur_pos <= 0;
            chart_id <= 0;
            seg <= "";
            state <= MENU;
            text[0] <=  "=======    Main  Menu    =======";
            text[1] <=  ">>> Score History               ";
            text[2] <=  "-----      Chart List      -----";
            text[3] <=  "    [0]  Free Play              ";
            text[4] <=  "    [1]  Tiny Stars             ";
            text[5] <=  "    [2]  Song 1                 ";
            text[6] <=  "    [3]  Song 2                 ";
            text[7] <=  "    [4]  Recorded Song          ";
            text[8] <=  "                                ";
            text[9] <=  "[^][v] Move Up / Down           ";
            text[10] <= "[<] Auto          [>] Play Chart";
        end
        else begin
            // Pointer actions
            text[1][0:3*8-1] <= (cur_pos == 0) ? ">>>" : "   ";
            text[3][0:3*8-1] <= (cur_pos == 1) ? ">>>" : "   ";
            text[4][0:3*8-1] <= (cur_pos == 2) ? ">>>" : "   ";
            text[5][0:3*8-1] <= (cur_pos == 3) ? ">>>" : "   ";
            text[6][0:3*8-1] <= (cur_pos == 4) ? ">>>" : "   ";
            text[7][0:3*8-1] <= (cur_pos == 5) ? ">>>" : "   ";
            
            case (cur_pos)
                0: begin
                    read_chart_id <= 0;
                    seg <= "HIS     ";
                end
                1: begin
                    read_chart_id <= 0;
                    seg <= "FREE    ";
                end
                2: begin
                    read_chart_id <= 1;
                    seg <= "SO    01";
                end
                3: begin
                    read_chart_id <= 2;
                    seg <= "SO    02";
                end
                4: begin
                    read_chart_id <= 3;
                    seg <= "SO    03";
                end
                5: begin
                    read_chart_id <= 4;
                    seg <= "SO    04";
                end
                default: begin
                    read_chart_id <= 5;
                    seg <= "SO    05";
                end
            endcase
            
            // Input key actions
            case (user_in.arrow_keys)
                 UP: begin
                     if (cur_pos == 0) cur_pos <= 5;
                     else cur_pos <= cur_pos - 1;
                 end
                 DOWN: begin
                     if (cur_pos == 5) cur_pos <= 1;
                     else cur_pos <= cur_pos + 1;
                 end
                 LEFT: begin
                     state <= PLAY;
                     auto_play <= 1'b1;
                 end
                 RIGHT: begin
                     if (cur_pos == 0) state <= HISTORY;
                     else begin
                         state <= PLAY;
                         auto_play <= 1'b0;
                     end
                 end
             endcase
        end
    end
endmodule